`timescale 1ns / 1ps

module NextState(N1, N2, N3, N4, N5, Floor1, Floor2, Floor3, Floor4, Floor5, A, B, C, D, Aplus, Bplus, Cplus, Dplus);
    input N1, N2, N3, N4, N5, Floor1, Floor2, Floor3, Floor4, Floor5, A, B, C, D;
    output Aplus, Bplus, Cplus, Dplus;
   
    assign Aplus = (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & ~A & B & ~C & ~D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & ~A & ~B & C & D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & ~A & B & ~C & D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & ~A & ~B & C & D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & ~A & B & ~C & D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & ~A & B & ~C & ~D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & ~A & B & ~C & D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & ~A & B & ~C & ~D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & ~A & ~B & C & D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & ~A & B & ~C & D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & ~A & B & ~C & ~D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & ~A & ~B & C & D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & ~B & ~C & D);
    assign Bplus = (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & B & ~C & D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & A & ~B & ~C) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & A & ~B & ~C) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & A & ~C & D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & A & ~B & ~C) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & A & ~C & D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~B & ~C & D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~B & ~C) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~C & D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~B & ~C & ~D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~C & D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & B & ~C & D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & A & ~B & ~C) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & ~A & B & ~C & ~D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & A & ~B & ~C) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & A & ~C & D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & A & ~B & ~C) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & A & ~C & D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~B & ~C & D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~B & ~C) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~C & D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~B & ~C & ~D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~C & D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & B & ~C & D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & A & ~B & ~C) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & ~A & B & ~C & ~D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & A & ~B & ~C) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & A & ~C & D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & A & ~B & ~C) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & A & ~C & D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~B & ~C & D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~B & ~C) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~C & D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~B & ~C & ~D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~C & D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & B & ~C & D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & A & ~B & ~C) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & ~A & B & ~C & ~D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & A & ~B & ~C) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & A & ~C & D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & A & ~B & ~C) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & A & ~C & D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~B & ~C) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~C & D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~B & ~C & ~D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~C & D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & B & ~C & D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & A & ~B & ~C) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & ~A & B & ~C & ~D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & A & ~B & ~C) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & A & ~C & D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & A & ~B & ~C) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & A & ~C & D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~B & ~C) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~C & D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~B & ~C) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~C & D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & ~A & B & ~C & ~D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & ~A & B & ~C & ~D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & ~A & B & ~C & ~D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & ~A & B & ~C & ~D) |  (N1 & ~N2 & ~N3 & ~N4 & N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & ~B & ~C & ~D) | (N1 & ~N2 & ~N3 & N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & ~B & ~C & ~D) | (N1 & ~N2 & N3 & ~N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & ~B & ~C & ~D) | (N1 & N2 & ~N3 & ~N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & ~B & ~C & ~D) | (~N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & ~A & B & ~C & D) | (~N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & ~A & B & ~C & ~D);
    assign Cplus = (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & ~A & B & C & D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & A & B & ~C & ~D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & ~A & B & C & D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & A & B & ~C & ~D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & ~A & B & C & D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & A & B & ~C & ~D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & ~B & ~C & D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & B & C & D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & B & ~C & ~D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & ~B & ~C & ~D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & B & C & D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & B & ~C & ~D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & ~A & B & C & D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & A & B & ~C & ~D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & ~A & B & C & D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & A & B & ~C & ~D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & ~A & B & C & D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & A & B & ~C & ~D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & ~B & ~C & D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & B & C & D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & B & ~C & ~D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & ~B & ~C & ~D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & B & C & D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & B & ~C & ~D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & ~A & B & C & D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & A & B & ~C & ~D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & ~A & B & C & D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & A & B & ~C & ~D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & ~A & C & D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & A & B & ~C & ~D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & ~B & ~C & D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & B & C & D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & B & ~C & ~D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & ~B & ~C & ~D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & B & C & D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & B & ~C & ~D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & ~A & B & C & D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & A & B & ~C & ~D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & ~A & B & C & D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & A & B & ~C & ~D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & ~A & C & D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & A & B & ~C & ~D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & B & C & D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & B & ~C & ~D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & ~B & ~C & ~D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & B & C & D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & B & ~C & ~D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & ~A & B & C & D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & A & B & ~C & ~D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & ~A & B & C & D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & A & B & ~C & ~D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & ~A & C & D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & A & B & ~C & ~D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & ~B & ~C & D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & B & C & D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & B & ~C & ~D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & B & C & D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & B & ~C & ~D) |  (N1 & ~N2 & ~N3 & ~N4 & N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & ~B & ~C & ~D) | (N1 & ~N2 & ~N3 & N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & ~B & ~C & ~D) | (N1 & ~N2 & N3 & ~N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & ~B & ~C & ~D) | (N1 & N2 & ~N3 & ~N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & ~B & ~C & ~D) |  (~N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & ~A & ~B & C & D);
    assign Dplus = (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & ~A & B & D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & ~A & B & C) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & A & ~B & C & D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & ~A & B & ~D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & ~A & B & C) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & A & ~B & C & D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & ~A & B & C) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & A & ~B & C & D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & ~B & ~C & D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & B & C) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~B & C & D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & B & C) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~B & C & D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & ~A & B & D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & ~A & B & C) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & A & ~B & C & D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & ~A & B & C) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & A & ~B & C & D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & ~A & B & C) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & A & ~B & C & D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & ~B & ~C & D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & B & C) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~B & C & D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & B & C) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~B & C & D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & ~A & B & D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & ~A & B & C) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & A & ~B & C & D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & ~A & B & C) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & A & ~B & C & D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & ~A & B & C) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & ~B & C & D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & ~B & ~C & D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & B & C) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~B & C & D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & B & C) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~B & C & D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & ~A & B & D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & ~A & B & C) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & A & ~B & C & D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & ~A & B & C) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & A & ~B & C & D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & ~A & B & C) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & ~B & C & D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & ~B & ~C & D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & B & C) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~B & C & D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & B & C) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~B & C & D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & ~A & B & D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & ~A & B & C) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & A & ~B & C & D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & ~A & B & C) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & A & ~B & C & D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & ~A & B & C) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & ~B & C & D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & B & C) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~B & C & D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & B & C) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~B & C & D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & A & ~B & ~C & D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & A & ~B & ~C & D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & A & ~B & ~C & D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~B & ~C & D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~B & ~C & D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & A & ~B & ~C & D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & A & ~B & ~C & D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & A & ~B & ~C & D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~B & ~C & D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~B & ~C & D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & A & ~B & ~C & D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & A & ~B & ~C & D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & A & ~B & ~C & D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~B & ~C & D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~B & ~C & D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & A & ~B & ~C & D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & A & ~B & ~C & D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & A & ~B & ~C & D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~B & ~C & D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~B & ~C & D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & A & ~B & ~C & D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & A & ~B & ~C & D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & A & ~B & ~C & D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~B & ~C & D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & ~B & ~C & D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & A & B & ~C & ~D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & A & B & ~C & ~D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & A & B & ~C & ~D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & B & ~C & ~D) | (~N1 & ~N2 & ~N3 & ~N4 & N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & B & ~C & ~D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & A & B & ~C & ~D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & A & B & ~C & ~D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & A & B & ~C & ~D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & B & ~C & ~D) | (~N1 & ~N2 & ~N3 & N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & B & ~C & ~D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & A & B & ~C & ~D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & A & B & ~C & ~D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & A & B & ~C & ~D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & B & ~C & ~D) | (~N1 & ~N2 & N3 & ~N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & B & ~C & ~D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & A & B & ~C & ~D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & A & B & ~C & ~D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & A & B & ~C & ~D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & B & ~C & ~D) | (~N1 & N2 & ~N3 & ~N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & B & ~C & ~D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & A & B & ~C & ~D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & Floor4 & ~Floor5 & A & B & ~C & ~D) | (N1 & ~N2 & ~N3 & ~N4 & ~N5 & Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & A & B & ~C & ~D) | (~N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & ~Floor3 & ~Floor4 & Floor5 & ~A & B & ~C & D) | (~N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & ~Floor2 & Floor3 & ~Floor4 & ~Floor5 & ~A & ~B & C & D) | (~N1 & ~N2 & ~N3 & ~N4 & ~N5 & ~Floor1 & Floor2 & ~Floor3 & ~Floor4 & ~Floor5 & ~A & ~B & ~C & D);
endmodule